package sim_file_pkg;
	`include "trans_arbi.sv"
	`include "mem_trans.sv"
	`include "drv1_arbi.sv"
	`include "drv2_arbi.sv"
	`include "gen_arbi.sv"
	`include "agent_arbi.sv"
	`include "arbi_monitor.sv"
	`include "score_arbi.sv"
	`include "arbi_env.sv"
endpackage : sim_file_pkg
